`timescale 1ns / 1ps
`default_nettype none
//////////////////////////////////////////////////////////////////////////////////
// 
// Module Name:    UART_Clock 
// Description: 
//
//////////////////////////////////////////////////////////////////////////////////
module UART_Clock(uclk);
	//port definitions
	output reg uclk;
	
	always #5209 uclk = ~uclk;

endmodule
`default_nettype wire
